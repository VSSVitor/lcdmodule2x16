library verilog;
use verilog.vl_types.all;
entity lcd_example_vlg_vec_tst is
end lcd_example_vlg_vec_tst;
